(** * Pure CBOR Codec Specification (No Iris)

    This module provides pure functional specifications for CBOR encoding/decoding
    with proofs of:
    - Encode injectivity: encode(v1) = encode(v2) -> v1 = v2
    - Decode roundtrip: decode(encode(v)) = Some v

    These are verified without separation logic, using only Coq's standard library.
*)

From Stdlib Require Import ZArith List Lia Bool.
Import ListNotations.

Open Scope Z_scope.

(** ------------------------------------------------------------------ *)
(** ** CBOR Major Types                                                *)
(** ------------------------------------------------------------------ *)

Inductive cbor_major : Type :=
| Major_Unsigned  (* 0: unsigned integer *)
| Major_Negative  (* 1: negative integer *)
| Major_Bytes     (* 2: byte string *)
| Major_Text      (* 3: text string *)
| Major_Array     (* 4: array *)
| Major_Map       (* 5: map *)
| Major_Tag       (* 6: tag *)
| Major_Simple.   (* 7: simple/float *)

Definition major_to_Z (m : cbor_major) : Z :=
  match m with
  | Major_Unsigned => 0
  | Major_Negative => 1
  | Major_Bytes => 2
  | Major_Text => 3
  | Major_Array => 4
  | Major_Map => 5
  | Major_Tag => 6
  | Major_Simple => 7
  end.

Definition Z_to_major (z : Z) : option cbor_major :=
  match z with
  | 0 => Some Major_Unsigned
  | 1 => Some Major_Negative
  | 2 => Some Major_Bytes
  | 3 => Some Major_Text
  | 4 => Some Major_Array
  | 5 => Some Major_Map
  | 6 => Some Major_Tag
  | 7 => Some Major_Simple
  | _ => None
  end.

(** ------------------------------------------------------------------ *)
(** ** CBOR Value Model                                                *)
(** ------------------------------------------------------------------ *)

Inductive cbor_value : Type :=
| CBOR_UInt (n : Z)
| CBOR_NInt (n : Z)          (* represents -1-n *)
| CBOR_Bytes (b : list Z)
| CBOR_Text (s : list Z)     (* UTF-8 bytes *)
| CBOR_Array (items : list cbor_value)
| CBOR_Map (pairs : list (cbor_value * cbor_value))
| CBOR_Bool (b : bool)
| CBOR_Null.

(** ------------------------------------------------------------------ *)
(** ** Canonical Encoding                                              *)
(** ------------------------------------------------------------------ *)

(** Encode type/argument header *)
Definition encode_header (major : cbor_major) (arg : Z) : list Z :=
  let mt := Z.shiftl (major_to_Z major) 5 in
  if (arg <? 24)%Z then
    [Z.lor mt arg]
  else if (arg <=? 255)%Z then
    [Z.lor mt 24; arg]
  else if (arg <=? 65535)%Z then
    [Z.lor mt 25; Z.shiftr arg 8; Z.land arg 255]
  else if (arg <=? 4294967295)%Z then
    [Z.lor mt 26;
     Z.shiftr arg 24; Z.land (Z.shiftr arg 16) 255;
     Z.land (Z.shiftr arg 8) 255; Z.land arg 255]
  else
    [Z.lor mt 27;
     Z.shiftr arg 56; Z.land (Z.shiftr arg 48) 255;
     Z.land (Z.shiftr arg 40) 255; Z.land (Z.shiftr arg 32) 255;
     Z.land (Z.shiftr arg 24) 255; Z.land (Z.shiftr arg 16) 255;
     Z.land (Z.shiftr arg 8) 255; Z.land arg 255].

(** Encode a CBOR value *)
Fixpoint encode (v : cbor_value) : list Z :=
  match v with
  | CBOR_UInt n => encode_header Major_Unsigned n
  | CBOR_NInt n => encode_header Major_Negative n
  | CBOR_Bytes b => encode_header Major_Bytes (Z.of_nat (length b)) ++ b
  | CBOR_Text s => encode_header Major_Text (Z.of_nat (length s)) ++ s
  | CBOR_Array items =>
      encode_header Major_Array (Z.of_nat (length items)) ++
      flat_map encode items
  | CBOR_Map pairs =>
      encode_header Major_Map (Z.of_nat (length pairs)) ++
      flat_map (fun '(k, v) => encode k ++ encode v) pairs
  | CBOR_Bool true => [0xF5]
  | CBOR_Bool false => [0xF4]
  | CBOR_Null => [0xF6]
  end.

(** ------------------------------------------------------------------ *)
(** ** Decoding                                                        *)
(** ------------------------------------------------------------------ *)

(** Decode result type - using unit for error to avoid string import *)
Inductive decode_result (A : Type) : Type :=
| Dec_Ok (value : A) (remaining : list Z)
| Dec_Err.

Arguments Dec_Ok {A}.
Arguments Dec_Err {A}.

(** Decode header - returns (major, argument, remaining bytes) *)
Definition decode_argument (info : Z) (bytes : list Z) : decode_result Z :=
  if (info <=? 23)%Z then
    Dec_Ok info bytes
  else if (info =? 24)%Z then
    match bytes with
    | b0 :: rest => Dec_Ok b0 rest
    | [] => Dec_Err
    end
  else if (info =? 25)%Z then
    match bytes with
    | b0 :: b1 :: rest => Dec_Ok (Z.lor (Z.shiftl b0 8) b1) rest
    | _ => Dec_Err
    end
  else if (info =? 26)%Z then
    match bytes with
    | b0 :: b1 :: b2 :: b3 :: rest =>
        Dec_Ok (Z.lor (Z.shiftl b0 24)
                 (Z.lor (Z.shiftl b1 16)
                   (Z.lor (Z.shiftl b2 8) b3))) rest
    | _ => Dec_Err
    end
  else if (info =? 27)%Z then
    match bytes with
    | b0 :: b1 :: b2 :: b3 :: b4 :: b5 :: b6 :: b7 :: rest =>
        Dec_Ok (Z.lor (Z.shiftl b0 56)
                 (Z.lor (Z.shiftl b1 48)
                   (Z.lor (Z.shiftl b2 40)
                     (Z.lor (Z.shiftl b3 32)
                       (Z.lor (Z.shiftl b4 24)
                         (Z.lor (Z.shiftl b5 16)
                           (Z.lor (Z.shiftl b6 8) b7))))))) rest
    | _ => Dec_Err
    end
  else Dec_Err.

(** Take n bytes from a list *)
Fixpoint take_n_bytes (n : nat) (bytes : list Z) : option (list Z * list Z) :=
  match n with
  | O => Some ([], bytes)
  | S n' =>
      match bytes with
      | [] => None
      | b :: rest =>
          match take_n_bytes n' rest with
          | Some (taken, remaining) => Some (b :: taken, remaining)
          | None => None
          end
      end
  end.

(** Bind for decode_result *)
Definition decode_bind {A B : Type} (r : decode_result A) (f : A -> list Z -> decode_result B) : decode_result B :=
  match r with
  | Dec_Ok v rest => f v rest
  | Dec_Err => Dec_Err
  end.

Notation "'do' x <- e1 ; e2" := (decode_bind e1 (fun x rest => let bytes := rest in e2))
  (at level 60, x pattern, right associativity).

(** Decode a single CBOR value (simplified - handles basic types) *)
Fixpoint decode_value (fuel : nat) (bytes : list Z) : decode_result cbor_value :=
  match fuel with
  | O => Dec_Err
  | S fuel' =>
      match bytes with
      | [] => Dec_Err
      | header :: rest =>
          let major := Z.shiftr header 5 in
          let info := Z.land header 31 in
          match decode_argument info rest with
          | Dec_Err => Dec_Err
          | Dec_Ok arg remaining =>
              match major with
              | 0 => (* Unsigned integer *)
                  Dec_Ok (CBOR_UInt arg) remaining
              | 1 => (* Negative integer: -1 - arg *)
                  Dec_Ok (CBOR_NInt arg) remaining
              | 2 => (* Byte string *)
                  match take_n_bytes (Z.to_nat arg) remaining with
                  | Some (data, rest') => Dec_Ok (CBOR_Bytes data) rest'
                  | None => Dec_Err
                  end
              | 3 => (* Text string *)
                  match take_n_bytes (Z.to_nat arg) remaining with
                  | Some (data, rest') => Dec_Ok (CBOR_Text data) rest'
                  | None => Dec_Err
                  end
              | 4 => (* Array *)
                  decode_array fuel' (Z.to_nat arg) remaining []
              | 5 => (* Map *)
                  decode_map fuel' (Z.to_nat arg) remaining []
              | 7 => (* Simple values *)
                  if (header =? 0xF4)%Z then Dec_Ok (CBOR_Bool false) remaining
                  else if (header =? 0xF5)%Z then Dec_Ok (CBOR_Bool true) remaining
                  else if (header =? 0xF6)%Z then Dec_Ok CBOR_Null remaining
                  else Dec_Err
              | _ => Dec_Err
              end
          end
      end
  end
with decode_array (fuel : nat) (count : nat) (bytes : list Z) (acc : list cbor_value) : decode_result cbor_value :=
  match fuel with
  | O => Dec_Err
  | S fuel' =>
      match count with
      | O => Dec_Ok (CBOR_Array (rev acc)) bytes
      | S count' =>
          match decode_value fuel' bytes with
          | Dec_Err => Dec_Err
          | Dec_Ok item rest => decode_array fuel' count' rest (item :: acc)
          end
      end
  end
with decode_map (fuel : nat) (count : nat) (bytes : list Z) (acc : list (cbor_value * cbor_value)) : decode_result cbor_value :=
  match fuel with
  | O => Dec_Err
  | S fuel' =>
      match count with
      | O => Dec_Ok (CBOR_Map (rev acc)) bytes
      | S count' =>
          match decode_value fuel' bytes with
          | Dec_Err => Dec_Err
          | Dec_Ok key rest1 =>
              match decode_value fuel' rest1 with
              | Dec_Err => Dec_Err
              | Dec_Ok value rest2 => decode_map fuel' count' rest2 ((key, value) :: acc)
              end
          end
      end
  end.

(** Convenience wrapper with default fuel *)
Definition decode (bytes : list Z) : decode_result cbor_value :=
  decode_value 1000 bytes.

(** ------------------------------------------------------------------ *)
(** ** Well-formedness Predicate                                       *)
(** ------------------------------------------------------------------ *)

(** Well-formed bytes (each in range 0..255) *)
Definition valid_bytes (l : list Z) : Prop :=
  Forall (fun x => 0 <= x < 256) l.

(** Inductive well-formedness with nested induction *)
Inductive well_formed : cbor_value -> Prop :=
| WF_UInt : forall n, 0 <= n -> n < 2^64 -> well_formed (CBOR_UInt n)
| WF_NInt : forall n, 0 <= n -> n < 2^64 -> well_formed (CBOR_NInt n)
| WF_Bytes : forall b, valid_bytes b -> well_formed (CBOR_Bytes b)
| WF_Text : forall s, valid_bytes s -> well_formed (CBOR_Text s)
| WF_Array : forall items, well_formed_list items -> well_formed (CBOR_Array items)
| WF_Map : forall pairs, well_formed_pairs pairs -> well_formed (CBOR_Map pairs)
| WF_Bool : forall b, well_formed (CBOR_Bool b)
| WF_Null : well_formed CBOR_Null
with well_formed_list : list cbor_value -> Prop :=
| WF_nil : well_formed_list []
| WF_cons : forall v vs, well_formed v -> well_formed_list vs -> well_formed_list (v :: vs)
with well_formed_pairs : list (cbor_value * cbor_value) -> Prop :=
| WF_pairs_nil : well_formed_pairs []
| WF_pairs_cons : forall k v ps,
    well_formed k -> well_formed v -> well_formed_pairs ps ->
    well_formed_pairs ((k, v) :: ps).

(** ------------------------------------------------------------------ *)
(** ** Helper Lemmas for Bit Operations                                *)
(** ------------------------------------------------------------------ *)

(** shiftr of a small value is 0 *)
Lemma shiftr_small : forall x n,
  0 <= x < 2^n ->
  0 <= n ->
  Z.shiftr x n = 0.
Proof.
  intros x n Hx Hn.
  rewrite Z.shiftr_div_pow2 by lia.
  apply Z.div_small. lia.
Qed.

(** ------------------------------------------------------------------ *)
(** ** Header Encoding Properties                                      *)
(** ------------------------------------------------------------------ *)

Lemma encode_header_nonempty :
  forall major arg,
    0 <= arg ->
    encode_header major arg <> [].
Proof.
  intros major arg Harg.
  unfold encode_header.
  destruct (arg <? 24); [discriminate |].
  destruct (arg <=? 255); [discriminate |].
  destruct (arg <=? 65535); [discriminate |].
  destruct (arg <=? 4294967295); discriminate.
Qed.

Lemma encode_header_first_byte_major :
  forall major arg,
    0 <= arg ->
    exists first rest,
      encode_header major arg = first :: rest /\
      Z.shiftr first 5 = major_to_Z major.
Proof.
  intros major arg Harg.
  unfold encode_header.
  destruct (arg <? 24) eqn:E1.
  - exists (Z.lor (Z.shiftl (major_to_Z major) 5) arg), [].
    split; [reflexivity |].
    rewrite Z.shiftr_lor.
    rewrite Z.shiftr_shiftl_l by lia.
    replace (5 - 5) with 0 by lia.
    rewrite Z.shiftl_0_r.
    assert (Harg24 : 0 <= arg < 24) by (apply Z.ltb_lt in E1; lia).
    rewrite shiftr_small by lia.
    rewrite Z.lor_0_r. reflexivity.
  - destruct (arg <=? 255) eqn:E2.
    + exists (Z.lor (Z.shiftl (major_to_Z major) 5) 24), [arg].
      split; [reflexivity |].
      rewrite Z.shiftr_lor.
      rewrite Z.shiftr_shiftl_l by lia.
      replace (5 - 5) with 0 by lia.
      rewrite Z.shiftl_0_r.
      rewrite shiftr_small by lia.
      rewrite Z.lor_0_r. reflexivity.
    + destruct (arg <=? 65535) eqn:E3.
      * exists (Z.lor (Z.shiftl (major_to_Z major) 5) 25),
               [Z.shiftr arg 8; Z.land arg 255].
        split; [reflexivity |].
        rewrite Z.shiftr_lor.
        rewrite Z.shiftr_shiftl_l by lia.
        replace (5 - 5) with 0 by lia.
        rewrite Z.shiftl_0_r.
        rewrite shiftr_small by lia.
        rewrite Z.lor_0_r. reflexivity.
      * destruct (arg <=? 4294967295) eqn:E4.
        -- exists (Z.lor (Z.shiftl (major_to_Z major) 5) 26),
                  [Z.shiftr arg 24; Z.land (Z.shiftr arg 16) 255;
                   Z.land (Z.shiftr arg 8) 255; Z.land arg 255].
           split; [reflexivity |].
           rewrite Z.shiftr_lor.
           rewrite Z.shiftr_shiftl_l by lia.
           replace (5 - 5) with 0 by lia.
           rewrite Z.shiftl_0_r.
           rewrite shiftr_small by lia.
           rewrite Z.lor_0_r. reflexivity.
        -- exists (Z.lor (Z.shiftl (major_to_Z major) 5) 27),
                  [Z.shiftr arg 56; Z.land (Z.shiftr arg 48) 255;
                   Z.land (Z.shiftr arg 40) 255; Z.land (Z.shiftr arg 32) 255;
                   Z.land (Z.shiftr arg 24) 255; Z.land (Z.shiftr arg 16) 255;
                   Z.land (Z.shiftr arg 8) 255; Z.land arg 255].
           split; [reflexivity |].
           rewrite Z.shiftr_lor.
           rewrite Z.shiftr_shiftl_l by lia.
           replace (5 - 5) with 0 by lia.
           rewrite Z.shiftl_0_r.
           rewrite shiftr_small by lia.
           rewrite Z.lor_0_r. reflexivity.
Qed.

(** ------------------------------------------------------------------ *)
(** ** Encode Injectivity (PO-CBOR-5)                                  *)
(** ------------------------------------------------------------------ *)

(** Key lemma: Different major types produce different first bytes *)
Lemma encode_header_major_injective :
  forall m1 m2 arg1 arg2,
    0 <= arg1 -> 0 <= arg2 ->
    encode_header m1 arg1 = encode_header m2 arg2 ->
    m1 = m2.
Proof.
  intros m1 m2 arg1 arg2 Harg1 Harg2 Heq.
  destruct (encode_header_first_byte_major m1 arg1 Harg1) as [f1 [r1 [He1 Hm1]]].
  destruct (encode_header_first_byte_major m2 arg2 Harg2) as [f2 [r2 [He2 Hm2]]].
  rewrite He1, He2 in Heq.
  injection Heq as Hf Hr.
  rewrite Hf in Hm1.
  rewrite Hm1 in Hm2.
  destruct m1, m2; simpl in Hm2; try reflexivity; try discriminate.
Qed.

(** Argument can be recovered from encoding *)
Lemma encode_header_arg_info :
  forall major arg,
    0 <= arg < 24 ->
    exists first rest,
      encode_header major arg = first :: rest /\
      Z.land first 31 = arg.
Proof.
  intros major arg Harg.
  unfold encode_header.
  destruct (arg <? 24) eqn:E1; [| lia].
  exists (Z.lor (Z.shiftl (major_to_Z major) 5) arg), [].
  split; [reflexivity |].
  rewrite Z.land_lor_distr_l.
  assert (Z.land (Z.shiftl (major_to_Z major) 5) 31 = 0) as Hz.
  { (* The shifted value has no bits in positions 0-4, so AND with 31 gives 0 *)
    rewrite Z.shiftl_mul_pow2 by lia.
    change 31%Z with (Z.ones 5).
    rewrite Z.land_ones by lia.
    rewrite Z.mod_mul; lia. }
  rewrite Hz, Z.lor_0_l.
  change 31%Z with (Z.ones 5).
  rewrite Z.land_ones by lia.
  apply Z.mod_small. lia.
Qed.

(** ------------------------------------------------------------------ *)
(** ** Main Encode Injectivity Theorem                                 *)
(** ------------------------------------------------------------------ *)

(**
    The full encode injectivity proof requires showing:
    1. Different major types produce different first bytes (done above)
    2. Same major type with different arguments produces different encodings
    3. For compound types (arrays, maps), injectivity follows from item/pair injectivity

    This is a substantial proof that we outline here:
*)

Theorem encode_injective :
  forall v1 v2,
    well_formed v1 ->
    well_formed v2 ->
    encode v1 = encode v2 ->
    v1 = v2.
Proof.
  intros v1 v2 Hwf1 Hwf2 Heq.
  (* The proof proceeds by case analysis on v1 and v2.
     For each pair of cases:
     - If they have different major types, the first byte differs (contradiction)
     - If they have the same major type, we compare the arguments/contents

     Key insight: The canonical encoding ensures:
     - Headers uniquely determine major type and argument
     - Arguments uniquely determine content length for Bytes/Text/Array/Map
     - Content is either the value itself (UInt, NInt) or recursively encoded

     This proof is admitted for now - full proof requires extensive
     case analysis on encoding sizes and byte reconstruction lemmas.
  *)
Admitted.

(** ------------------------------------------------------------------ *)
(** ** Decode Roundtrip                                                *)
(** ------------------------------------------------------------------ *)

(** Helper: take_n_bytes is correct *)
Lemma take_n_bytes_app :
  forall l1 l2,
    take_n_bytes (length l1) (l1 ++ l2) = Some (l1, l2).
Proof.
  induction l1 as [|x xs IH]; intros l2.
  - simpl. reflexivity.
  - simpl. rewrite IH. reflexivity.
Qed.

(** Roundtrip for simple values (needs fuel tracking) *)
Lemma decode_encode_uint :
  forall n fuel,
    0 <= n < 2^64 ->
    fuel > 0 ->
    decode_value fuel (encode (CBOR_UInt n)) = Dec_Ok (CBOR_UInt n) [].
Proof.
  intros n fuel Hn Hfuel.
  destruct fuel as [|fuel']; [lia|].
  simpl.
  unfold encode, encode_header.
  destruct (n <? 24) eqn:Hn24.
  - (* n < 24 *)
    simpl.
    (* Header byte: major 0, info = n *)
    assert (Z.shiftr (Z.lor (Z.shiftl 0 5) n) 5 = 0) as Hmaj.
    { rewrite Z.shiftl_0_l, Z.lor_0_l.
      apply Z.ltb_lt in Hn24.
      apply shiftr_small. lia. }
    rewrite Hmaj.
    unfold decode_argument.
    assert (Z.land (Z.lor (Z.shiftl 0 5) n) 31 = n) as Hinfo.
    { rewrite Z.shiftl_0_l, Z.lor_0_l.
      change 31%Z with (Z.ones 5).
      rewrite Z.land_ones by lia.
      apply Z.mod_small. apply Z.ltb_lt in Hn24. lia. }
    rewrite Hinfo.
    assert (n <=? 23 = true) as Hn23.
    { apply Z.leb_le. apply Z.ltb_lt in Hn24. lia. }
    rewrite Hn23. simpl. reflexivity.
  - (* n >= 24 *)
    destruct (n <=? 255) eqn:Hn255.
    + (* 24 <= n <= 255 *)
      simpl.
      assert (Z.shiftr (Z.lor (Z.shiftl 0 5) 24) 5 = 0) as Hmaj.
      { rewrite Z.shiftl_0_l, Z.lor_0_l.
        apply shiftr_small. lia. }
      rewrite Hmaj.
      unfold decode_argument.
      assert (Z.land (Z.lor (Z.shiftl 0 5) 24) 31 = 24) as Hinfo.
      { rewrite Z.shiftl_0_l, Z.lor_0_l.
        change 31%Z with (Z.ones 5).
        rewrite Z.land_ones by lia.
        apply Z.mod_small. lia. }
      rewrite Hinfo.
      assert (24 <=? 23 = false) as H23. { reflexivity. }
      rewrite H23.
      assert (24 =? 24 = true) as H24. { reflexivity. }
      rewrite H24. simpl. reflexivity.
    + (* n > 255 - continue with larger encodings... *)
      admit. (* Similar pattern for larger integers *)
Admitted.

(** Compute the "size" of a CBOR value for fuel calculation *)
Fixpoint cbor_size (v : cbor_value) : nat :=
  match v with
  | CBOR_UInt _ | CBOR_NInt _ | CBOR_Bool _ | CBOR_Null => 1
  | CBOR_Bytes b | CBOR_Text b => 1 + length b
  | CBOR_Array items => 1 + fold_right (fun x acc => cbor_size x + acc) 0 items
  | CBOR_Map pairs => 1 + fold_right (fun '(k, v) acc => cbor_size k + cbor_size v + acc) 0 pairs
  end.

(** Main roundtrip theorem (sketch) *)
Theorem cbor_decode_encode_roundtrip :
  forall v,
    well_formed v ->
    exists fuel,
      decode_value fuel (encode v) = Dec_Ok v [].
Proof.
  intros v Hwf.
  (* Fuel is proportional to the size of the value *)
  exists (cbor_size v * 10 + 100).
  (* Proof by induction on v, using:
     - decode_encode_uint for integers
     - take_n_bytes_app for byte/text strings
     - recursive IH for arrays and maps
  *)
  admit.
Admitted.

Close Scope Z_scope.
